��
l��F� j�P.�M�.�}q (X   protocol_versionqM�X   little_endianq�X
   type_sizesq}q(X   shortqKX   intqKX   longqKuu.�ccollections
OrderedDict
q )Rq(X   linear.weightqctorch._utils
_rebuild_tensor_v2
q((X   storageqctorch
FloatStorage
qX   77766944qX   cpuqM�NtqQK K
M�q	MK�q
�h )RqtqRqX   linear.biasqh((hhX   77006880qhK
NtqQK K
�qK�q�h )RqtqRqu}qX	   _metadataqh )Rq(X    q}qX   versionqKsX   linearq}qhKsusb.�]q (X   77006880qX   77766944qe.
       �Y����?!��?�X뿎�F?�'A���M@����$�㿠      $8A<=�	=x�<*N��,����o�<(	�<���G|���|�<
A�<��<��<"4�<�Y�<�ɍ�<�7<S�ʼ�}�<2��<���"J�Ω)�N0M�@�=�����$S�<�v�<�<�;ʣ��p�M<�;��`�O�<>k<��;< s0��w<O�<0�2�/m�>H�>�4�>L���V?V�>Zo�>m��L�<�Ƽ\�Q<�� ;��I�H�;���/^=��j����<���8P>�q;>�4������h�>�<讙�Ҷ�if�8?"���c�_���z=�s���	��)�����_�@�r���R��76����� #[9��c<�9����nꆼ���a|���?�+�����<@a=jo��T�.�Ĳ>���2��=��=�)Ż6��;��=��.����XJ>4��i,���>�n���>�{ɾp�D��a=�����=�q�5;ͽ������D����=x�.��2&>E	�.@�=�Ƕ�j�=��!����=�>���==ŋ(;��<��<�V���-�=��<Y��ѻ�>�ξ(<<�u~<Rm��;�6����Ǜ>�>��Ġ>�ٽ�[��[t<�1�=)]!��q�� =��_<ؠ�<�z&<:���<s�<-�f�����#=h|ɽ�+��
���;������=�6�<�&ӾZӾ���=7�;�m�:��ּe�=�� ��q&�ݓ_:�ϝ�G��=��Ҽc�4<��<뙼�d=�<mO���O�=�=!���_�Խ�!M����򌽸��K��:*����+ݾ"�m=9��=�>=`�z=7���d�=1B<<!2�=��}��R< �,=J����Cg�=��;8�=���I�»�t̽8��=70y��:�=~��e<�?"fC��bL=~X2?Y����6&��U�g̻��k�	 �</_��wJ� ��=`�y�a9�=?d��/�=B=`�<�g�d^=Q�(=�\>�5˺k�<�u�m9	����⯫<���<��>�Mu���1<وͼ�%��\����~=S>u<ӝ�=�wP:��%��|�=<P=��k���<i�<(��<��A=R� ={F�+C��=�E>=>�Q�UcܾP�)�.^�c�F�[I?%徽��>��9>S/(��1���Շ���K=c�J��=��L7T9�A'=E+d=$�`=��'=9��=�!��3Q=)�z��|�=��<�=<��5=1A�$�ʻp�l<�[�?�~��ǫ=jGC��%����<!�=2UG=�}6��}�D=�@��ga9=��w�u���A܈����=�.ʽf��<��q>��B<�=�6������5 �Q=��-�Qo��f8��ާ�U%B�@�A=���=�d<[μE�X= >p���<�}=ǭ=q���;X����<�..<�Y�+�����=x����=S<�j�<�g>�`��j���s�7�3<<V=���YJ?�'�>���.��<ܮI�k�;= 5��-�s=�*=��ּ�e�`$!<��+58�3f�nuF=���<�C��4�4��Ō=���=Iz���>_U��=@��`V�;n�����;I���Z[�����=��+=�	�=	n��H�=⠪��ł<�u�=��<"�@�׾/=ƒ�A�u;�ܼ��5���=7�=���;��=��C9�Pw�B0[��� r%<�ľ�w�	�+����2?>�:[<d��R �=^S<=��@=h��=�颽`��<�K��A#���O��Z��)�m�>�;��!�<��:�=�Z�<ƓU>��u=S��t�!<����&!�<��X��}���H�5�=�-�<{�&=U.=��=���.u|=W������]���=�_�m�<����n�<=ܷ�K�(=�����O��r��Q	�0�y�o,�?��;J����L���"=��=�K��=���<3	��X�s<}U5=�h����<Q����ϼ�F���`9=�kG=W����^��=w���=��j��&=�ڤ=o^��Iy?Dw�<f��<(\� >���=�*���-T<�+?�Ҁ�=��z=}?=;�<�ُ��C��eQ���<�����������|��Bѽ��;��-����=�ҟ�z >޸Ⱦ��1�8�Ҽ.�>Z����\<�矽Ke=EQG=�o�=C��D��Z^<Z��)�=Kt��h�<�&���<<����S�<.�����=��7=)+�=����t>$�K�<뻾�p���ʼ`��>��6�4�4z'>>��=�H��<f�,=}44�;e�=�<�L�=D�<eV��@�=☺����<��w=L R��.(=yG�m��<S�9�V��Gj�\a�<���4�R<@t�:�WU����>�r���B*���P=.4X=�iP�Ҙ�;̮I='� =Yӱ=�S�;��?��p�<�v=����!���d>��7�l����=�Ľ�Œ=������?�$������Jz�Q�Ծ:|�#��߇}�i�=��?�l�%=�V=�d];�\ܻx�	�(>����ʈ�<���<<�m=�x6�0�=�s=;���#>]��=�Z����>��/?@�ƺ"�<�|= ��<:D�K���N�=�̯���=.��'ˬ<Pک<~2F=.�`<׽g���=�&<sӎ����=w�ؽU�����;�%�
͘=@w=#�ݬ?�վ��W�z�ʼ*��<��KTɽ���>g$�=���O�;��=ceӺs�=�,%�J�>7�;���5<?�Y;�D����e=���=�m~�ɍ�;�t��U֋<�������=O[�f��<|$#<�?������V������+`Ҿ�/n�R�-������=�J����?>�J��qf�<��e�}��78�~b������H����l��#�Ͼ��׾α��;4�� ���=N�����U�UQ�P4�<@�<<��A�:�Q��+N�'V����b;Rƾ ���\l�P��y1[��z���`��^�����ի;M�[���P(�tX��ӄ =X�	���< ����K$��P��m����k��b<P{�<��Z�r��<1�@�	������2��e����.7��W�<uyͼgi`<*�<���F2�;:��A d�a��������< aκ�E�xEW<��Ѽ)B=~rռ�P< �Ǽ�¼�<r��< ����l�X� �"���ŻlȼF��H�����<���<ȳx<`��1m=P�Q;0���=��R��<`��;.:�<�l�<"Y�<�<<��=p�7<�;��Z<�p�<q�=���<������:B�;?� ���= �5<�$���E����)������Y'��o����<И;��<\\ɼ�J���Ż<|�@�0�d;�^@��V��f����;�	��6�����=��5=�᝾���>+(Խ�P�>� >��R>v���|��>���>q�c��g����HӼ U��£�<�s<�]��N��<��><ߌ>Q ���ϣ��/��=;����O���e����|NU=��=N�{��=�̽za=� ����=�Pk���5=K@=}��>�V義�G�-���pai<���:���պ�>@в��D>����/>��žR��>��=䪚=\��<�4���;t=���r�<�;�m���JY=��$�<֚(�Q+_=�I���ܿ�߮���z���O�<���=�N
>|Ē>rΡ>�>���F:���s���2�YaQ��o4�4���HVɼ�7=�aX<.�]�H�z<���X:;��<ͱ�=�����u>�s�H�
<�$��'� ����z���e=W�>T>���Z�>P��{=�q����c2�<��
�����\�ڼ9����A��Yy<��/������=��\;�ގ�=�j��N�^��sμ�j�<O)�ߠ����&����>w}�������4>��(����=O2�<�/޼�=��?�#c�;�*���<)����%�_`#��.�=�\=zF��|�̼��U�O��J�=���<B��<�]��*ܽ]�1�vr'>9D>'D�qN��QsS��
���*Z<<��е�<�/�;�s^�)�H������=>�<�<�ݎ����[�
=�@x=�����W4��Ѣ���'��:��,�Y��ͽk�,���
>�-�`n�=��?>Y �<s1;����:�;�1����v<��<I�=v�!=�C�����<I�����<w;�==��2��c�>Z?b���>-I`����:��a�#��׾�G$��)�{�.��ݫ>'g>���<w��=YZ��lp=�=�}=Kڌ;��&=1�D�==KDǽ[%�<�F�<-y�=�N�$: =���=��?n�ռ��G���>I�\�Z�K>���>��Ӻڽ'����!���c�ܑl:��ܼ��r=^
=	�= B�<nx�p��;��d�����>kJ��tP�>�;0���w>"}>i^=?�Ė��U �M�Ծ�2�=~ς>т"��{�=@�>v��}W�=	T�;-���<k=nS�=�R=��E����<�.2;��{��1��B�T<��k	?����"S&>b*�;J >H�̻ �@<�O��IᎽYr�=j*-����=��=j{�<�"�=H׽��ؼ�0=SZ�<��<cѫ<(�V=�%�<��漳}����%=h��|x_���s��̫����M��=�t�<LYͼ���~E=�<=d�?��>z�Y>�dǾK>�=|B���<rA��f;Ψ&<Ӊ�=��&=д�;F;�86�4�-��<-�=2�y�\�=�@�>(&`�j�>r?qS�h�ּX,<ܡ�=��]>'F�;���U�V��Ve>��=�ټ��H�ղ�� y=�gN=2��=(���s�=�c�xr�<'���D�j	���&������Ǿ���=��>��p�y�=@����=,�$�T�<>�(����-��]��=�tz��ͤ<�0��R:;d�5=I^(��ڻ<�*ؽ!�Ľ��M���=��=O��=G{�B� ?˵̾��=�j���M�<����郼�����=:�����e>_�<�IR<W^��kZ�<Wi9�
=裄=g=7��<#ka=&㑽�������=�܎����\`/>ͽ���_�=,Uf���=��=��<��9=�;�s��l2�*Xȹ�c�����������<Z�+�k9Ѽ@�Q�?��e��<��n<7@ �lõ=��<Oؽ1��=h$��8t���4��yq&>X�:�O����>＃=�=!�O=پ�=��=8�����=��>�zO��ϊ=-��<�����q.��'==&���UQ=���=7��@���M_�=.J��_|��(D>����2=���=61=��l>`5
<[���M��v;��b��=�
�����[�`�VCD<I4:��<���<0=�=P��Sg�<�cU<��b=��=le=�i6;>��sX�=�8��~>>(� A�>�y=��>�9�=MW˹��>;����#=�Ĕ=5�=�lʻ��<��=�s�?��
X<%�=�=?��<�J�<���=��ܼ�4���>����jW���m?Mb�=x�= 1C�M�J>?��=H'�e�<6�=�]�>���<p%�� IL=�g�<��9�d׶���V�0���l;��� G��=D��=t��<�>U�>��Ͼ�$%>��v��-#?=�j����< 꿸�8R;[��<��f��M�W<�@�{W�<ܝ�~=�����n��g�<��f<k���=�+=�s�<4�J=X��[=��[���&<��>�A��C����[>u��>�IݻJ/���<<Ө<`�?H����an��U����z=Q�����߻ٷ=ƍ)�v�q�4(+�w��<d���_�>�J/�K�>�R��=⽋��:=����hk�>WL�>�큼z��<�'�<��_�&yĽ���q^K�ã>9`d���3<��L=��D�0���=>��Ӽ��G��LV��M
���xA}�f��ە������w �͌�<�:~<��< _�;�e�<Ѝ��Hq�;#I�<+����a;͛����gT��I��=�$��(��S��!<��R��>�M���Խ,r���yԼB���a��S/������:����X��P� ;�	�;�Jy�]�< DF�x�;$O�<���<�7�<S�<�����̼^[��ѿ��V�����t������(�������*<IP=N)������м��W�l=�7D<�P��r��<ꤦ�Ќ����̻���<�9�q�=P��;z����x=�"<��p<�-<Gm=�ͨ<�y�<�=p%[��
=4}<�|�< :2��<B�\�<�1��I=�<��<Ű�w��`~�<0l������>�Zq��d=?T0�!W^�@?���=���\�<'J>��<S��>��!�Ϟ=��������٨<<�L�|���hz<P�;��Ź6{�<��; ��<2�r�=�_>~���*=�>(��=�	�=p��=L���Q�;���=dMA=�C=X�>�ǽ�=7>��>����z�>�I?c��=�U�: ԼCq߼��l�k��;�m�*.��&=��Լ���=C1��>�/S����==o�<�->��<���<�p=`FU=�9�hkA=�d��֛=D�~=�ξ��Q>�R�=��!�j8��Q�:a󜼛����x>������$= �b>� ׼�%�<��*=�M�=7����4=���*Ir=,�C���=/��;5L�<� 9LH�<��9�n���9���T<?u�@�Κ�r��.��<7/>�#=3\�>�;�3�<�0�<�"n<����yvm<�̶��:p<z��;e��<=����=��/�Ý	<Q:�����:v�<�ҋ��=��O����=�G��y����u�;p��=�Z�7V��&=
�<�.=D|�<܊^<C&A=N���=�;��漰=3�;2GK�?���};�9�f��N������tڽ�΃>��
��;�	�<��ϼ*�>�K>;�=0L9=���<"Jb�ҸG=��뻌e����2=u�s����<���<{���l�<�^�)sD<
vļ�&��lq�<�`g=�T&��3����J>��Ƚ�z�: ��';�>p�X�bړ� p�=��L��<�B<lx��o�E<Z�U=�zY��J�����;XZ����ںA�(�nJ'=���W9�<�Ԉ<U�$��}ʼ�I�=5�6�[;��%�5������Q�o���ё.��=�o(<2�=�~��]<� ���8�<���<�8%��(����w��4�:;�*=�T�<�BX�ne-<f͐���;��]����<��=����!Ͻ]�.>��&�|"��ˬ�V��>ҋ>o׽�9�=���=����3�<��)���S��J<U�.��M<�$�<�3���M;�*T=�#o;C��
9�;,=��d���3�	�U�>���-?+7�%2��p����<���u�<
�;=�=ׅ6��j�$�=������ھu��Ң��WT��̼!q�F�o�3-����!=p�v�EGT=2�<"�=N7E�y�5>�+~��^��Ɠ<R+[<BA���	S�tJS>j
4��۽�N�M�S�એ�?��<f�����˼d�Ƽ��ռV`μZ��@�XW�j�C<XA<������<�� �>�8=�>�?�>��c��a�<�a;��_��
%>�7��n�<��j���ؽ�=��E�n�8����<`ʮ�2�`< I�;#�v��N��+l<�5�'�<����;�<Y�»/׼e�E>���=�I�>}�>z|ּ�[.��)�x�*=���=��k������rA= r6;'3Ƽ���<�$m�<4�7�0�
��<�[���̻[V�� ]=��%�3%<&ix�����ă=���ѐ�<0�>눌?xY�<�-��/(>�D߽� k=SJP>���=џ}���<��Y=���Ji<�/�����;�Q<�߻��H<�/%��
G����<��0���I=͐�����1�>0��=^
��[�>����/��Xd�;�ō>u=.<��;S��<Ni=ۑ����Z<�X�;]��<�X<(2=�I�<�	���py<\ٴ=:p�;r��;�T���'S=q��<b��=<*P=!�q>���>�*�>H|���н���>,˵;�k[=�/�<�{=
r��t�<;�;2&=�9�<wA5<<�3=!r�:�!�<�%=b)<��[;�Һ-J�;[1"<@�N<���<1D�Ja>��)=v��?��X<�Zm�����'�=�׳<k�=���<Ȏ�=M�������}�T=ȥ�<�1~=�n<�Y<p�;$��:>g+=�%<%=k=�˓<x�=��=<p>D�X>�lg���/>�<9�ܤ�c��ԓ�Đ�<�]y��b�;��F=z(��e=@��<���<��7<�1�=�CM<�=�=�j=엺����^ڹ<�Ά�0�O=�=�q��w#m>�NT>��׽��Z��8`4>A
>_�x=Z�=�t=��]=>�=Z�<Mx<%�o=�u4<�P�<��e����;x��<*:��;�=�5;�ʟ=�H=�z8=�ҥ�y��=Њ�=J`��G�:�p��k�8=I�>�N�=����6���i���<!>�ND&=�	����<~U�:O!�<QM	=��t����<?GI=V�<4��=�9�K=������Y>�K��� �>]Z>r+�����?
�:� >z��=� =�#=B�j=���<<�,={�3=���<��;�<��><		�A4�<�<����~�Q=?��T�=H��;�R={5_��J">Nܑ=a%�\X�<�����U;Ī=4��=_>����<v��<���B<�%��$����<1�Q�"r�<�ڤ����<4Ag�Vl�<�Ɛ=Rx"=���<e��=8f�>���gd>�GϾp:;5ܼ>��<�Ď�"9O�cy�9ĥ����<�C��><@+�;����
�<�x=���^f�=8q�sM�=`=�Ƥ<p���ZE>Kv�;�����f?�ԇ>LR�>>Ȯ��=V��0ũ���ռ���ϕ����>�����R���m���=�?(�Mn�=�k����ػ� >H1��	>�2(:�"L�߫d=�RT�������Ծ�C��
�5�Zp�>J��<��<��< V;<@¿;��o�=�����ӽ=�Y��z\�e���&6��X��&�s�bŞ�0�� �S���S��럾B�|�P�弿�1�x{+�)���5��<`A�:�����;Ǿ��#=#���8�Q<����TX<���<
�ʼ�<)�d<�܅<�'w���ڻ����(Q�@g��5���	�kF<��<���6C����d�kf��p�<Α< �:P�3;��W�.C�<�=�7g<��<�s�<A��$�h<�`�<����8�<n���fn�<�<��<~��<0�i<�%B;,��:��<�=���<h+�;����Z�t�<  u<��=�\�<�:���<J���"o<��k<V͵<�%C;�F�,�2FI�擩�o��<��������ek��!|���Nf�	�<�,>�|�"��w�< �z;Տ케;��<��M<ҭ�<��мnM�<Бż�I�����<�
1�p�4�<'ؽ��N�Z���<�~�<�*�=>6*��!�>Ns���>W|�=ݠ�;�=���9�>��׾�&Խ��>��,��T ;�Q
=��Ѽs=��!�J�߽|S��ޒ��Q�=�';��{�2�}>Z�=i�> `�<9�>�V��]�=3C$<��=C�˺8Q�=JW�^Y#>H�c�D�O�p]ҿP�F������;P$�<`��:���<��<�U��񾽟��=��'>��
���=�oA<A̠=�	�;i�<�)=r��<�HK<�K=�'���H�<��<=��\�(�k��=𮾲p�>�~������!��ńƼ.值���;��=M�4>[�=`4��.5�=�����=�6����<\U<�l<�<�<��<p��:�Y����9<�ߵ�G��t�r<5��=�&���TN�:<���@�<R	�<Y++>��|>���=���;<=P �<c���U��<~��<@,=QcD<�
<��!=�(6��*d<���<�)1��Q2=�i̼Zք<��+=�+�#-4�o��=��辇�����\��,�L�>N_=�~>�|�=T�s=�*=ꦌ�X�G=W�O�V�~;�۱;��<�޼l!
=��<���<��<���I�<9�u<�]Ѽ���gQ<B,:�r��[����<yu��C=w��i >�:=�C<Á#=T�<k[���r�w��<��,;A�B< ��:K:�f/��P�<�c;>(=����g;��O;�D=������ʼD�_�a�<�T<<x�[:�D1�d	�>d����$>���μ�<��;;k�=��=�Ы�F㘼,&����;_�=Q�=���< �=P�<��<�=��C<�o6=��ż�>�hX�>�N��\�����*<Z�=��P�J@=]6��f�=EZ$=T�)��ố���퇼�N���
-��]�<��л+��<�S�;�8<�B<ἔ<��<����FV}���=D{����N=���萼pȽЂ���-�����>%>?��a��:������X������l
��늼LU�<�S5;��<���C˔<��
<e�d��\�<���#k�<���=n.=�$8c>�����<I��������V�<���W`~;�=<[q����9E�f����9@ED=,?�B}�<q�>��?=DM�;�<}*�F�<;�<.*�<n逽U�w�E2����0�>����6=2�,�&���,�b��B>׉2��C>S��徰�Zo�;�}�;7�f�o���W߻z@F<���<9<���g�<�vŻe&\<8��<aq���:���ֽ-8�=L��=�ړ�\$��͖˼P�����=����z>�4�=cnG�l���W伋b�;�k���<,"���2�<]|;�<�<8��;��W��_�;1��<�_��ܼb�<�t��m<7=����
�l�غ0��X����=6P�=1���_;��h=��H<-���s��밼�f%�R;�r�<E�T�mBY<��
;w=�<�r��=ͼ5H<�e=/��;�<%=m��=a�;==F���T�>��[�!=\�A>��>���=:��=��L�̷T��,ͼ�r��Q�<6�5���<�Z�j��=U����_�;%IQ�Hb:��=�B<_v�<�� ��8=9��2�8>69��_I�<�����<F�>����B8=�`�=�4P;�r�< ,�<�����Y������ �a�x�y���Q�),��j�=2��<sɿ���=�9�[=�p;��<�C���Ĵ������������P$�<��>M�=���;1,L=��0=Us��5E�<��=�[�5�ĝ��Z1f��6�����<�=�`�<�̈<6n<� ��<[,=�%�<Jު=/"=��v���k���S���׼F~%�ʧ�<Y����P=�W#<U��=�d;�L�u^�B�O���Q;.:�g�;��;�r;k�L<�	�<U+=��<�+p;ߙ	<*X�8S�����<�����`�3qA;c���j����+����4<�6>�v�=��=��r=Ϊ�<$) <E=��\�	cƻ)�8��l�<�V<'¶����<H
�<s{�<r���v�|="gQ=���<���=��{<f���p>P,�;�̧�	*:�y�0>-U=�B^=pƼ?ֺI:)<3�r<檻�L4"���Ż�{�<5���a�<�D�<��%=�}9��9�<<=J��$ɔ��+�;�*=��3������C>��=Wǽ}���`�<�m>�ڊ= Bq�6=~/�;k!";2(=P���ž<>���ٻ�_�F��<rr<u(+=�2�;
���V=���I��=Mո=��P��{�<��>�=���l
�<1��>(l7=���=�o=�=�0:=���<�Â��q�<8�<�K��U��=���#�=O�����d;�R=��<l;=�-=� ��xY=\��3���5�>�;���}�����?�>���>
o�=�Q��F�=��<6e�<���<���<�m_=���rB=��<��,:W�<�=�;<'�1���;qh�=s�I=%{>�fT�j/���L��F��t0<�Y�ģ���_��:��@>S��<h��=`U>��=���=��;4�=�v+=h'=��=�O=�<���=y>;>�xn��n�M<>ZF��"'�5+�� P��)�<pGA;�= �X�ɔ����ƾ�s�>غ�=�+">Ẁ=�%;���=���=�?��]�i=�E�=�Dm=%�=�ޟ=/(;K��^�>��4=1�;�7۽�=�����w<���<f� ����<��=�F<�H;:��<8����`��ݝ�h´Aƽ�m�i^#��
ٽSk*�����l��_(���e1��j6�ԯ��\�< t��y���=�N�<+� ��y��)�= ��;�E(;�<ƃ�<�٫;�E��n!<�_�<H:μuj
����L@<z��|�@1���纼��Ϻ�R�@O�<����Z(<tR<�o=x��3�;�M��A��@.�$Oj<Ӗ=}�<q�Խ�Ľ,	�m$�.�E��r��俾�k��4p�>�����߾ؽ;�zr�ՠ�uD����������y[D���;�ۖ��L�< W��w ���<�hF�fW���Z�"������oX��Gv�����F��4�ʿYK�>$$�P�>��<�Y-���
= ľc�<��ھ,Z���qb>�����/���<2q�<��#��=���N�i�B5��AԼ��>�I��8ƾv^>��߽'2ƽ��־]S;�Y�vl���8�=���Š�=Zhڽ�tl=��=̓��=�]���������<X��<�m<��y�žp�>w�"=IE���U>m�C�[r�;o13=�uG��EͼH=y{!�t��-�<A{c�)�a��ғ<'��=&�=�q>���=Q�z>�%=����yt�F	���<>k�����>y�s<�%�=���=6���8�`=�}W=�%�VYK<��=Z0'�fڴ</��<���o|�<���;|p.=Gq����1	��Ƈ�<�-g��=�h>�z�p��;�s�#}�װ7��c4=9>����t�|28�'=1$�$5����E��	�z���͒V��@��ۓ��b��A.�	8[��W�X�F�f!H=�=�أ=֥<\�Q�󢭼�#*�ŉ��J>�k�_�=�B[=��g<I]����<�"��͚�9�oB��vD���ȼ��n�{�&:;U�5��d�</�;�D�<�=��d=��0=�q���)>�e��뗾ߣ��;�?m�>Œ[>͎=pq��z�<�ռ`^�<>	��ҋ�<t�������W���m"�Gc��.N<��o���Ǽ�=(���E�H��i�?>��
jɽ �غak9��@�>�yB���ҽ���<�r0=��;������;�<ټ|=����G�=�������<`�:�U<�&ٻx,< I!�0`(= �=橡�����BK>�˄��R�;�a{��d�<<�T�r�<]���`�k�
�<�v�<���<S�����0:!�;<ȓټy-�u�<�X����<�¼*B<��4�<$L�<EŽ�z�=6S���Y��ZD��`�@<_����-=��S>YA�;GHt=&=b2Q����;��f=.�u=!�:�uޥ=����bc��+A=�^P=y��;��<jл�j������Ysn<���Z�ޞ)�q����ٸ���麃h��A�=Rt='=���=z�M=���=S7=��;gq�<�/=(Ƅ=�E*=�uj�$��;��=^�;�D<v�<�%<<#p�=:�<@}=�-i>)N��ʏ�/6��>��<�%=��f<eF^��lG=_R�~F��aW=�d�<+�X=��n=,� =�U= ���N7<��9=&��<��;��%=�z,�i�<��=�s켻ᶼ%H��?>Ue^>n�u���=���=��L��F>?>F��=]Ҳ<��{<Yh�<���;L.�<�R�<��=� �ü =�k�;̩0=�=%/�
H=+T�<��M;�Ӟ=/�~�z�=Z�>�$��ᐾݭ =�=��9?V���^=5Fi<19J=	70==��<DZ=ֽ�<Y<=��\��ѻ���;`�<TS=��?=����6�<)����d�
>q$=�p���a��|ب>S�c����< ң<��ž��_����08�Y>��X�<Eߥ=s�q<��]�����*B=�ͣ<�t�<[��<���<��=S$=�_7<
�U=��a=VI���=��=6��< ���m�>���< I<ŋ�>�7�xFT�/�<�0Q���u<�j9��y�<ə�� ��<�ü�T�<��<n2=�i=_�'=��H=�H�X����B<���<\n.=3�h�֚�<�б=�TB���ؾ`q�<X>����Q�9=>$D�u�d=���<��<O=��-�4}"<E�<wd#=�yF�+�<#�w=�hƼ�����(=��=�=W⍽���=�C=�p��Dr���G>���<%3��(���:�>��Լ��>	�N�L�?<t<���w�#�μ�Zg=�E��Pܻ|=Tx�Hؼ���+�G�̅j�q�G��b�=�����6�'%��^���(>�<l��<�N<vi�=y�꽼\>�����Z>������ý�^�<�|���<E���9�`��;O)��=�p�<%㸼X����R��
�;�T���n=�.y�ZjĽl���Y����m<����rqq>�P>�e���[�>�p�v]�q��=k5=Tԓ��%:�*��<�F��;}����<2�1�	c�<��I<B"�<t}�=߳j�r�?=~0)<��=���<���i�=�;���ӂܼE	���n�޹g�Ǚ=Xm�k��4+/�����' �'���W�tqּ�����<���;�D5�^�=����L�=w��=R��=�7>W{ľ�
?# ̼И��V��<~�ż8v���U��N�uus��ì<	�K=l��n�ƹ0J;���^&<TJ�;#��<N <�Di<-�<n�4�=��<�=��l�1������>�0��30:?��<��ټ�$�;�x=���{������=��>&d1;���~�h<���jp�=VP�Z<c�＀R���<J��ޗ`��!�=24���Tl=<-> s/>��9�p��?������<�h�<^ =���@��:]�?����`��<�n���#��$B=	K���TR����;hV�<9s�<��_:c�"�ƒ=¬�S�=��<�r!��k�w>�	� ⓽�33�غ_<��i<L����=*1Ľ�x^=�>vgI>G�ξn�=*����0������}���rT-��Z��8ֺ;W������Q��"�:�XPU���ʽE�=V�>�h�<�dy������<����Ҽ(��;�C�:2?(�9��5��z��d��K��(������i���C�뾝���P�������˽M���.8�A���T��U��@$}:J�<����];^D�<�	�<���<���;��`�F�	��.μ�����=:�<�+ܼ��<
y��(��;�-��(��;����<Rh_�X�<D��\h5<X0传����p�(;&���ȡ;��ἅC�>��< �|<,���!=p���`�����<@��:��*;@;����p�ἔ�d˄�����̳�<&./��qԼ7���^��<���끻dx˻pjg;�!=�<'����<LM���Fc�a��9���N��e��@�Ӽ���������wC��4=��{����C��H�=�\�v>���=��=D�5>aw�v�>�=��gb���W�nV����_�=�u�;Ў�<���=��H?����D�꾙�>6�U���p>����O]�=�s���q=FF=��%���<��P=[��<�w6=��i=tM�=����z��=/4t>>�Z>�'�<&�<jQ�<qg�d�>����H�����k=�4�=������<�R&<\�<ʤ�<B ¼�Y�<��<7�Z<�U�<�=�m=�w9�DR�=�;��<�Z]>c�<�T�B>e澘�S����"�>u�ʾ�
�;jy+��Q�=;��<�<��<�p�<α����:�+;̭�xc�<㾕<S��uf��u.=&�:A��<��<z�_���=�>�+�d<*��<�>3��k7>���=}�<B�-<B��t�<]䊹rk>�X�/=�1 ���G<�Y!<󕅼��;��B<�7=��w<�Ɗ�+Z�<�$4<�`�=L��=h!<���<�%O�`M�>���_m���o��|�;n����я=9cw���e<�<�ϕ<IB���Y�<\�4��<S6����=�<s�f<:"<��=��c<���<|�0>�E;65>�MH< �E�F?�T�s�B���m!2=>�<�Y�Ȼϧ�;b��<F<�� <�w�:�r�LB�f��<����AW���㺽�=��1;��;�K=cb>��M=K�p=��<:>�<��<;�q�>���ɇ�2�	��q=��^�ge<��b�u9��|7=4X:f��<��޺��/��T�'І<����������c=�@=�)=���=�'>WX�=w?��i�<�z��.<�n���K�=h�=��p���=a�T=�:=��=�4�<G�=�l<�X�<{Ɔ<U
�ȏ�����S.��ɑf�^]*={�軧�Y=��T>Ⴈ<��=Ȉ��`�;X���	��<X���(>��%��Y=|��$@�;�<��:�6�\<\Z�<�A=���;����E7	�t	��3�(�_�ɼ�.\��o��\����V<�W�>�5>�ʋ=f�
>t1n<叽y����ފ>�qx��<E({=�=&k�
�:k.=���<��</H�<��׻ѫ�<����U�+9)��I���-6�%��ؖ������}�
�T�>�S?M� �e��ʀ�~����n���j=�>y�޽� 
=�XϺ^�x;����<-=O	�<N�,��[ܼg�	����|��;}�=��{<끵����<>&���'��J�`��>����'>�[k9�[�<��
>~o'=�^��F$=�.Ż�a�<}�u� �>=*g�:X<�;A�<:��<(!�er���t��8tk�p�W�0z!<Ö�;'�\=Y(�eM�>M)�`��,m����#>��t�廔=���L=�o����=�4!<�_��Z��<Ck��X<t#�;1Hƻd~�����c{<����(j=8K�<�&:��E<��ʽ�==s#>���=�������I��{����,�G'�=ȝ[�R6t=q�6�L+x���P;��K����;�mR��ê<mF=:|��`hܻɛ�ٴ5;�ϼ߲�:�<��R��=�黒ُ���J=I�A��`��`�9��w�?������=9l�=�4 ��G�=�����@��T	����)����D���D�����U;�=�.�<(��<�<�|��T�=�w�8�,=��}=���R=ύD�j��<Sp�B۾�R=>��=�Y[=��C=�cO� 1W��]��~<���	i��`;r��;�r�<�m\:�Z�<��b�=[�p<�m��2�=R%c=���;,b �8I%>a3k;4�K<E�>�S �ϳ�=�f�<щ�=�Hz<�O�<�;�;Q.�<,�����<���;��.��f�<���j�E����;AF�9=pv=E����:�<�>��>Aj�����<�	)=2�="�">�ּ��'=Nu�<�Ԑ�Y�=f��<^�H:cL�<���q=�/<�U���=�S�<�ņ;&HU=�+��.U���c=YP�=�<U�D�g>F������=�Ս��S⼧,s�:��#��=z>2=z��#�<�"d<�Y<2_<�="��<�˶<p>2=�1�<0ƺL�5=�j���g����8=e2=��%=d��=��Oo�={�(��>�����<�7<�X>h��<,��=��m�¨�<BE�<�ݼD�=[`��:�<���<OI< ��<�]�<�m=��3;��>=ܠ[=]�o<�>=FX�0z:>Qn=4�ż�>S����,��$�i�>�mL>���=˩�=R�=w�����Q=�3�$q=�6;���<�P;�3'=���G`=lr(����H� =�ʋ=2�c<��	�'�>c���g��>���>`?N<�a(<Dk<y��9��<�1��D0=�=.��:痍:n&�<ۑ�;�=9����;=���<�#=?I\���e=��=[���qVL=��$�X�=� ��p�>:�����0�T;L,ȼ%��J6�<�B[>���>����,�=@@
>B/N����=J<�,�\�=,[�=Ѽ���=�q�;��=ެF=y�h>ݓ���B=&��>�Cg��`?��<��:�<B.�<�c�xQ
<`�A��������X�˾�*��%�B��1�;X��$$>&� =*�>X�����C>���=,>=3�r<&=��>A��=�q�u[b�ݔ��j�`��Pc���������<�v�<��ȐŻ��)��[P:�)�8��t��=�[�=8����:�<�#�V2ͼ�C��W���۽)�N�_�C�ux����\���E.����<0��;�I�\�@<�9�:H2�xa���d��t���(;U��� �@�@y��.<?
	=��E<�N<` <:��<H����<�[=��*<ECļ�M޼���<@I�;�>�<�=��
=*�]��%�;�=���x�˼Jv����ռp�->�P���Ap>�V!���34u�䋃=�o�={���/O=��<�>W�=��>d�>�n>�7�<�<ٴ�l$�e��1N=����������<=?s$F>*������X+�<s�=���=B�!>�%>�==9 d;W��=w'$��=U��=���=�t_=b.>G�>"�<�F�>�}������|�;�M�;&Ǜ<��f�]��8=�>�ɽ�½KW�>�>{1=��>�1=�6�=b	����R=Q��<�I=Be<��;5k4<��3=�$
;G�;=;�=�Σ=�G>n����?���<��=��<<6�����ﾾ��<��I>y���n�=�;E�!�I��<�2)������w����%�ڳ��:�< �[<
7������G<�)=��;aW�=����@���r�V�$?�ϻ�Plo<Ϸ*�Nib�5�=u�v����= �v^�=�}���a�=������;xT��BW=��d�(f��l����љ<�}�<�<�|�y=���d��=!��=�a򼤶^>ƙ�>�|Ѽ6#�<D��=�'���z=-e�=;Cm�J�=tAE����6���#��<��;�X��WcM���<�Q3���+<F�d�����㼃�=�O�+=�"�=�%�����=~Ɵ�_v�>��L��1�:��hy�����=�>e>��4�:}�=�����w�<��;Fd���6�~����K<�e5�dKK�^i��,���6c�����=òƽ�����L�>�@/�7�P=*.H>�h����<�3���K)���������w�=3��$$��7�:�7�:\���ar.��D=�x������^�ʥ�<�����֋�����o���ߡ=7{ؽ��N�f7=>�:�=[�վc�=\�R<s֙���=���>�����0�=�̠�u����ۼȲ��#݄��;��a:;v�+��6��G�Ƚ̺)�c����=�;�]=)w���%<����;w��*�e��xi<���<�Y�����C ���'�7'=6����8c=�"��;��8����O�<3kd�U�~� �;��
U9�u׼��콐�*�I����-μҏQ�4�=��v�4(��*P��:�؎
<�=;�H�U�A=��L>'��Sg=eI���7=��żG���fd;�<#�3��x��<-��{]>�r=�jK�_0�=�,����=4vi�xR!�g�<=�>�����@)��M�{�$��0�����U�<���<�p=C�e=Z<�ڗ=��C:��<�y�;ףE��!m�h}#=�^��}�ѽ%��U�չ=Ib�=G�>��-=s���C��/�=��z���|<�B��:�=`��=��= ?�m�6�s��[�<��t����<7<}�ٻ�s<���R���N���ƸF=2e=�Y}=��=�b�=�<l�=�V��,<� R;���<����&�������I�=G�<�����<B=>�0=6�}=ߖ���:�$��t\�:�=`���<�-�;D�<h3�;��޻�<�Q >�B>�2�=����n*�<�2ڼ��������[��Q�ǽ;��;Wn=�{�<�QJ��[=r�����-=9#�;�D=�U뼀Z�;O-)��X�;ɷ¼�L�<94<=��*���=yMY�f��=vx��{�a��[�;�+0�p����4��tt�>I�3=w�n=��9=��:$"w=�2�;�w�=��e:��Y<"���{��9_�3<F���F<�;�<lzW�I9,=��1����i؈=���=a.�=�����[<�;4ؼ;�Z��4ݾ�>ӛN��������=,n<	�=_�=����2
�<�V=�ټ�j�<E��;.G��Y�<N�-=wFa<��L=J�/=)���&y�=�,�o0��P��;H^<�b<�}n>��=������<z� >UK�V�=�P�;C��xڸ=���<C����=DeB�,��<$�<t('9"c�<=���&	="XW;~�[>j��	6������
��ǈ�l����f=�F=w��<c���!�<ȡ�<�?=�&�=^[T<�-�<�@b=��I=6�;���<�;�O�<�n<^��<�a�=���=s������;���[�,;j�A�*�<B�/��=ȯ=�̃=p�y��ڀ=v#I�w�=�{�=E����=�������=�=<sx=�*<�	= F���=s~q=�2&��b��w�<�W#>��A=����zw꼞
��=��jD��x���f�Gͺ��.<�==U�'=����=V{=��Z=Ì=W <=?=ĝ<;l[=w�#�f�5=�齽��@>� p=�>��'>]��<�ƻw����L�Fl8��<ٻ�U׾hu	�ߊ���>��4����<l��=����n=�8=Жd��H�=J�����x=��@��� =�7�;�W
>)��7�C����ɍ���D�>���)�;�=�G���9�Q��<�x!��n+���Խ�f⼖�=h"��__<��<�?߼�ҳ=XV/���= 5O���1=��=k(�<G����\>y�ξ����}�?��q <�I��7�<�1�����h&{< }n�������<�:��-+-���p�x�������a|?=�m8��g��<<:�=3	��S#>P���Ѹ�>�����Ⱦ��3���<a�= d4�>�<����������P; �2<�tڼ���?9���@~�4���#0�(�>'|&>�c���̾g��2�������@�3_���/�P����<kc�\g����]<`+���7�\<X��U뺌���ӛ;���<�L�;x��;z��<x�ۻ2��;�����	 ��w �M�a� ����c�0�;w�<ES���n�<��m<y���'�:h��; 0�8<�<2��<ϳ�;�<�:C;TFz����<G�5���x����@�<�Ui:@>�:kr����B��<��<r��<���<*��� >��:_����<��$����<��ʼ4�N<�X�<�������<�"*<%�
�\hڼ PӺ������D��<�qF�@ܓ;�^��7�<W�<JF��t�< �F�@Q�;S�<�S��Ф1����< ͒<F��:�<�+�<�EѺ$~޻@�|<��ͼ8�c<��&<d����+{<�G!<�T���2n��!�;���M������(I��Eѽ��ٽx?���������� �Z������U�<�8;X�T<��;^��#w��`a���<L��<87:���������<��W����<�=z��qO���û�+(</L�e���a׫��$���Ug�$��t����Q=�7���?W��fR��E��.R����'O�B^�<��Ҽ�O��Л<�5ۼf%�qL;9���:�(�T�����;˼�҄����`C����Ⱦ�þ�ؾ�]���Ϗ���,����W
��;�aj�.�� ��;h�;n/��`��:^��v���;E�S?[�V?z#��ٍs��H��F�<����=DN�=k�R���?��#<�va���y��m"����$���>�i;�댻�=S�<�a�<ހ��<:��,=��<���;<?d��v��J?��a�Zd=�~;=�6 >I`��^���U=]�<|@�;0i�wOL=�X���j<1�ؽ����*�k[9=(�	���<�hW��dF�Py�<������������>���3�=y�I=������=V�.='�2<�U�=J-�<�+<�k<�J4�Owp<О�<�x:о�<������=j	�<�L"��R<�O[�"z�����W��;Ϸ�>oX>��;>��x=oHS��G�=��=�qJ���0=Ye=��)<V��<z�	=��&=3�=b��<q�'=tX�� �S=	�==�,�:���=Ҫ��ͬP=�S�m���M�	�>,՟=v{�=�i�<^��< ���_�=n��=�j�<r=�<� S=>j=��!��V=�
3=���< ,���M=�8;�f<��;���;W�3=(�ƽ��9�Қ���B?�CF=�Ԅ>�ď=1r�=_�v=eԆ=<ʀ=��{��&�<���;���F��;��=� �;=+�=!H�<:B<_��=��<��=޺�;�x�<�S<ґ�<7�>�ߨ=t�����4?\����>��>1�=IO�=2�;I��=}�=E���W+=�E�A�+<�YE�2�=R��<��=��k=SO�9�<�;�8=�N�<�;=�C=�h"�(I�~�`>oa�=v�?Fv9=�C�^?�>��(<q�U=2�8=����'�	=���6s	==X�=V��<c�=D<(�=:"
=~5/=�Q={�=ǐ�#q�=���C>��Ž�]+<Q2ܾ��	��;�?ǂ�=s;�>2��=��=dkV=�e3�� Z=z��=��D��m���=��v�|Ӽ�C�:��Z=ӝ<=��*=��|=(��<exR�z"l�lA�<�M >/���3u� ��<'�?I�=I��=���>���=��=gW�<�=�覼��X���-�f�C<�<N���L�������;��<����^��.��f�=V�=J��:�'��j�>��=5�<��:��<q`O����>����ȩ=���=�ք�yt�M��<5R��ɺ���-��U�'�,�Ѻ0���@=��(=�@P=k��=�CK=_��*%=t}�= }�k��:���6�����Ԇ���F�8{�>�ѼR.<���<!,�;v$��搼��ۻ�B�;�΁�����
<��B=����=�<�8�Zl�<PL��_?�=��=�:�wy�<m料��?�p�e�n���X����<�=揁�h;ټ��X=���Ǿ��$��9½j�U;ܬV=�}��ȹ<)�<|�<�'�<	Vh=�[�;L�#=��9�	� =?10����'r�mi�V��<x����<A�/=�Q3=��F=p���Ѓ�;(2��J<�����¼�|<�~��/�<��<;9�;ܖr<��D�ڭ�*s=2~ƽ���=�h۽��i=�b=���>����aV�>��|=�@~>vK��a����L�=�*���f=����O߼�� =Cc�P^��v|=uf�<�I\�W�<�,�I�'=��<-�W���P=Ý��DH<jV-�9�3���)?)���N��<�>S�?��>��>w� �nS�=Z۰��յ�˪������H=9ǰ<sZ5�+��<�������?\�'���F�<��=�6�;��w�F$��P�>��^�]Q��`� �^��<���C?�X۾�=��Jټe���똽cc�</�����;��k�^A�<�W��w�<O=�^PƼooP�����"�R�=�S���;_��(e�=��=�$B����6�<���Q��<�����Rf���@>���=Т���(��c=M����v��d��;����\��5(�H��<h��;o��;�zǽ\C�5�[���)<�Ҽ���[OY>{�*��<p��; �C�t"�R%�NW�=����"<=
Y=;	h��hF=�����<}��Z�2=f1�:�@�m��<�Q$���>_1��W�u=�����������
?t��f�4��=<��=��ʾ�U`�NT)>D���7�?=��n= �6�Ƽ���������h�Ƽc�!��˂���� �L���#��ŽQ���5��=�XɽAt�>Ca�=�d��%贼pq;�m���=�[�=�ؐ�1��=[��<M�	=6��<v�n�
<�p�<@J^�[Ď=_Ϻ����<�a�;���<U�P���L=lR�=C�A�W0���k���k���C�����;�-�9&f3��mY�� >� �=꣊=2�e����<�d�</f=�=H�?=�z?=i��;��B=�t���<����X�=qI�S��<�2�=�;/=|vo�v�r����dﭻ@^��z��Ǆ	=�B�n�kш<=��0�=�$,>�x�<O�z=��=q.�<t��;���='�<=�}�=�Л=Iw�=�k�=��>|�;��0=3<�>*E�Z��ി����>=Ei��7�<`Rk� ��:�u�=ۼ>0�=�ރ�㰂>`Y�k�=���<n ��>�={G>ݰ�=��K<G	]>���M>��q��>�9K��3M?P-/<$��󭚼H)i<h�<<8+��;S<l���̺Ǽ��<JD���0<ni�� lƺ��;4 <���@�l���<�^y<�>ۼ��<�.<<��<n�R�������������2�h�J< &�8��; �Z9����̼�<V��<��=�>�q�=���l�;kD=�Y �h�����m�<-�;[]��J<��iH���
<������]ռ�������<���<��B��e��M=8F<0��<������<�j.�؁�-\=0#�'�̽�{��s����q�':�ė���/�XM4���Y�=�/>��T��G��+��˼���g;�?��C�ϼc���4d�6�"�<�ӽ�a�!=guY����Pk�/:�=�x�=p�V����=33�����=�$��v:1=�B�	�<�ET=�`K��1��J�=x��<f%�>�9����^>~nо�V�<�ۗ�9Z=�d&>L}���&�8�꽯�����Q<�I8=H/;G�D=cg5��=�-��~�=6):��={�<�L�<N��<��<�l:<�s�<r��/=>��<�"W>�*��#< P�9*�,�[����>�J�_��<O�b=�.��A=�	�c�=ŗ<�Ծ<L5�<< Ձ<�=��9k��< �%���b<�U��5<��J�<
��=Z��^\�<�����0����� ?�[n
=P�r<��<�|<��<��;�CQ��B9=ʯ��ȭ޹�8�<@ې;i�6<]cS��C=��;�_�;�w�ԙ�<�]=�=>�W�J�ͽ��<zP��l�,��=W�;���;>�	Os=�����:�J�[�u� �kK��R��<���<+��&�<caa;=+<�G�<a�A=�B�<a^�jQ=D~�=�gG����c싾o3��4*H>HS�=n�f<��`=<ظ<�Q��̑<�I�<���;�e"<���<�?���ҫ�wζ<ᥙ�'ު:Y��<㋅<X���Y�<���;�� >��=9=��H>l��Od�� _��)dg<�����X���J	=c�¼�n[=p�:�D�W��<󺼱�$<��;�涼�!�&ם<��̺��B<K��<E�<h�M=f,�؇>�� >@XԾ���<�6��D:��ʳ�����=�!<�C%=��N<g�.;^ <���<$�<���<��[<�kϻ&9N�Ñ��q��T�<{�=�3�� �o<��<·�;�Q<����ކ�<���=ǳ<u�^:����}�:��Y3=Qz<��C=�M=�)=K�=��?����<s1��ʰ�<��?=�����o����B*���Ƽ$��;�~���Pj=��<�R�=nǔ<���>1sF�|�������ʾ�%M>Y
=�Ҝ=L�.s?<����-<ja�<ɹ���[�<��<F�<���<�H�;��=�^�B"F=O�<�?\=#�a<+��<�7>�>r�A �=|a���f<�|��+о�y_="9����_�U�'�{K;=1Du<qsv<�	��R�<ʝi:K=z	�;P��<��J<��v��IS<#O�<�?2=����d�= 
�=K�ܼR��=ş�<t�(>�4ҽ�����<�L>B�.���=/�J=��ҽ������_<�2H<�n�<���<�R�<���;��ض_8�<0^<)���ȼzk=Qj�� ��V�a�{�F>/�>e)�\:z��h�<&��;r�2�C��=����~^F��u<v-�����<��I#����$<ă<-ۦ<}�q��򟺺�ȼa��<�-�<�ډ��@$����;�c�R
�;���<����=�B��ؼP�f�F��<Wm�=k�6��T/<�s<��	�8&�;n�R:^�*;���<qG
= G1=L�<<��:��<��=@�*���K��,[��b׼�$�$B�=�׽S>i�}mѻ���*��=��>h�>V�Ƚ\����*�<M=�<G�<��ǻ;�<�l�<L;��:�%0�xKA=���s����<5�ļ'�,=fG�<c�<�8>����6��Jм�����k<9	�������(��<���<��H�p<>F�9ǭ�<���<gTI<Ǩ5<BuغZ�<.cy��X�����:<[� �<��ܻ6�;$љ;B��{d>�P�۬��[p<��Q��;l�%g>���;쀇=�d<��k<�<�iZ<��x<g��:��
;�t�:�hi�鴅�e��:�G<�<ծ��v��<��!���L=]�p=��q�kՒ��g�r��H��<�R7�(�����u=���<ŭ���i<�� =tf<zp��7<M���^:Nj�<#n����;�0;L�:�C�ީ�;a�
=�=�=�F;�ܞ=�֡<��F=��{�м��嶽	�<�8�� ���.��<�2��C��<r�=A����=�9��{;
<�껪!Y<
�<d唻9�3<㪤<�<�;���<d���<0[=g��=Nk'�����2搾1�<-3n�Q3�*ư���>:=�^d=<�i�;Nn��b<�$;yϖ<��::><Gڻc%�<�E�s��<�Z�<�[y�0�;ǛT<�;<`�; ��=�I�=y`��>v�<�8@;�1�KϚ��	7���=Ô��Ny���%�<GQ=H�J+<'&��<�7=aĽ;d��<F)=�B<_��<��D=|���V�+=�?<�kB>V^�;����Ӿ�}�< ��<�
<�����W9���张�#�Z�#;���<�B;��<��%=8��<6��<��>;ް_�&�1=��Ѽ�VT=`OM=#�<��;�=^������FA�T�����������?��<�ۼ�2R�ޜ��C�=�Ֆ�1�0=����J=���&*�<��f;�X<s0�<2A=�ɸy=���<�<�=���<�I�<��/_Ľ&�"�-����Ѽ�I=��<�v<��a���ɻ�����t	�4"�����">v׼Q���7�=�&'=p婼�NX=e�`��m�<�+�n�+=e�t�&��S�$>�V8>��8>�
�'΃�}�=�
ʻ���:� =��;*#ʼh��*����
J��&[��.`9�mO�.��!�'���I�; ��'C�<�X��1F���h�#�ʼ��"����u�\�S�<:����,;Pڼ�>��6��<�Ȱ<�� <�vػ��ɖ�\fռ� ʼ��ռ\]μ�}� )�OO��>���>=���<0)�<��t=]<0�i<|[�<�����qL<Л�<8��V�<:��<�<����PŃ;b�<�w��N�<�)
�T�o<8:ͼ�X仠���!l���F��j�@t�;Ȯ�� ����-�� �a�`K��l]�����	�<����l��j�<2��<���<�'�<���#�̼*jx������D��n�<�Լ	 <w��<#�˼X�<��X��TO���f����Fˠ�^>���B\�z2R��I'�k6��h��<|Wo�{V=.�p��<��� ���|���˦94#��8z������f�<��*<q�g��$�����&w��X¾G�վ�,*�6D��ڢ�\�+>��
�t2���T"���8���&<]�<՝ܼ��b< �<�E�@�:�U���<��=��ý�}3�����R�����(�=#h}�)1��ͅ;�,=�
/�;Ь��� ��:=ۛ~��ޝ>�b6�.j���p��̫�<�j#�z&�@O��@o���R��U��y�N�K��T�@$��Ti�<ȪR���=,t�����=
�︹�!=a3���/=�2����'��$u�ṏ��h���(�7�P����3��k,��c��<����ȼ��,����8��d=�����<������C=��>=:����=���<N�@<�=j�޺3�-=��=�Њ<*g�<T���4�<][J��d=mc$��4>L����Q�J�^��돾;�Ľ�.�=�W����F�tp;a��(���a����;�6<[�< =���;;=��(=�\�<QS�<�qz;g@+=�{�;`��;G��<H�-�ӵ�<Mc���Ӿ<�:��Dj���
�����=��>D�ü�ܼ�2=]�;t����;�ʇ�+��=0M�:�<��s�1!n<�W����ì|=�6�P����8��� >��E�a'��͈�i�ͦ��|o/>Z%��e ��Zy=}��<��;+��<�J<;�<�<!W�<�;�;ʸ4=�݂�+o�<9�;�]���H�<:$7���=�<��b�<�z[��\��� �R�1���½٠+�=l��=v��&<�L6<�	B<4�m<�1���>�;_WK�xɰ�te]< ����
F7U^����\;DY�<�a'���<iS���$x<5w�ӉK>�F�r��̖�G80�1dK�f�d��Z�+=���9`�9=�[>=C9�<��~=��&<��b=Ֆữ8D<结<��<n��<'�<�x��?w�=�)��rx�=[�T�,;rׯ���>�T+�<&<�U�c�>#�=�x=8��<�=;m<�<�f�<�H�;�E=B �U�<F��<A�=87�<���;�'=�&=�k;m��=��.<z�g>n>���Kɾ�����W缰BO;��@�]�=��?��(�=�{���B��bm6=,t=g�;���<w��:�u��s��<���<�5�<�d=Aw1<C��<�.�<K��<���<�߸��D׽ܲ�=i�L�e�>j�5���?��ֈ��d���>nn)=5��<���<!i�ԏ���$;)�<����J��̳<1��<�T�:�=�2=o
=Td<��<�_]����<*�N��`H�!2/=O�>��{�+���¼��
��n+>�B��1��<<8=��<�,<����t��<<=���>��:'*	�?�<Rby�h�<����}�;3v�<�d��˩-=���<wa��:�Ｚ�>��j���;�Gj����=Y8�튉=�����?;��/��'=���j��<-Q<�W9͕�<e�X���I�˷=�b�<�<�Z�Oy~<��I�(*=�	�<ڬ����<�3�p>š��у<��[�\�ս<wd=p۽ێ=�����L�<�<q�V;�v;>����<f[<�q�k	=ն�<��0�;j��iO���x�����;����2pg=x	��sJ=n�j�Ґ��74>|���w>lt����:����H� =��׺f\�������V=�^=�r�[j�9�<Y��;��<� <\�M�/gE�%�<�=Q�w=��ҽ��/�[8n�]����"�P�<�Z���1���=��F�$g�i�6<�;����:���8�Ӽ��
���=�W������IӼNz��M�ּ:���(=)9j=H�$=s3ؽᩌ<EoD��O��Vd���jP������Xc��$_�pV���4=�ij�0df��cb<��I�|�޼�A�{�~�
Y�;Z��������;W%�<`� ����᳕��`�ƈ�=1^!=�(�=���>T#�h�<,���q<*FI�C�"<'���>��%=��g<Gj��2�<��Q�6�y�T<9���1�������>���̼�v:�P�<�qS<�B>#���\��
2>�Uܽ��A� P6<(�v<S��<�e��S
C=���>_*1�G�|��(j<&�<U��>�e=��ɻf��<s�W����<t*��C����F�<���:��l�AAF��½���<�d<>1�e>$㖽9
X���?���Ҽ��弱zྎX�>sV�5¼�8����<b��<��]X�b���J��o�ۻ�{�<(d�;/n���V��V1�p�=��i;�ԧ=�$�=k����>�������p�b<@�:�<�<�VȾu��@�~>5��=�o=��O=�,<T�Ȼg�;z�B<^�ɼO?/� �b�a��;d@W�*��:���<.�	=۪Y=p�E�T��=�y;>s���L0g>�樾"��<a��9c;;P>$g��+*1�
DS>�6����=Fq=R�)8��<=TT��*<3��;�J�=��8�H
=|ĥ<�U�=u��;��=�->2ʍ�]O�=�N���H?�Ε��َ�8y��hS��<��,>�6�>��$�=KG->�=|��=0 �=�C�=�R=�J]=rY�=���=���=(Ɓ=v�s=��=���=p
E=?Y=��>n?tG�<ʿ�<���<`�	<�I���˻@	�<���#���5=�(>F�-�=s��Ѩ�� �r=I���^�=5�v��� >sh���0!>ZB�R�r>�]�4\�=�8�Zhܼ���E��TJ�